.title KiCad schematic
.include "C:/AE/LMR23625C/_models/GRM1885C1H220JA01_DC0V_25degC.mod"
.include "C:/AE/LMR23625C/_models/GRM188C71E225KE11_DC0V_25degC.mod"
.include "C:/AE/LMR23625C/_models/GRM188R71C474KA88_DC0V_25degC.mod"
.include "C:/AE/LMR23625C/_models/GRM219R71E105KA88_DC0V_25degC.mod"
.include "C:/AE/LMR23625C/_models/GRM21BR71H224KA01_DC0V_25degC.mod"
.include "C:/AE/LMR23625C/_models/GRM32ER61C476ME15_DC0V_25degC.mod"
.include "C:/AE/LMR23625C/_models/GRM32ER71H475KA88_DC0V_25degC.mod"
.include "C:/AE/LMR23625C/_models/LHMI_5030_74437336022_2u2.lib"
.include "C:/AE/LMR23625C/_models/LMR23625C_TRANS.LIB"
XU7 /SW /VOUT LHMI_5030_74437336022_2u2
R2 /FB 0 {RFBB}
R1 /FBM /FB {RFBM}
XU4 /FB /FBM GRM1885C1H220JA01_DC0V_25degC
XU5 /VOUT 0 GRM32ER61C476ME15_DC0V_25degC
XU10 /VOUT 0 GRM219R71E105KA88_DC0V_25degC
R6 /VOUT /FBM {RFBT}
I1 /VOUT 0 {ILOAD}
XU3 /VCC 0 GRM188C71E225KE11_DC0V_25degC
XU1 0 /BOOT /EN /FB 0 0 /SW /VCC /VIN LMR23625C_TRANS
R4 /EN 0 {RENB}
R3 /VIN /EN {RENT}
XU6 /BOOT /SW GRM188R71C474KA88_DC0V_25degC
V1 /VIN 0 {VSOURCE}
XU2 /VIN 0 GRM32ER71H475KA88_DC0V_25degC
XU8 /VIN 0 GRM32ER71H475KA88_DC0V_25degC
XU9 /VIN 0 GRM21BR71H224KA01_DC0V_25degC
.end
